module multiplicacion(a,b);
	input logic a;
	output logic b;
endmodule
