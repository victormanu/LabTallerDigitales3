<<<<<<< HEAD
module ALU(in,out);
	input logic in;
	input logic out;

endmodule 