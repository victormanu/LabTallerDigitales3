module ALU();

	always @(*)begin
		
	end

endmodule 