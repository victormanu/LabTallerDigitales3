module ALU(in,out);
	input logic in;
	input logic out;
	
	always @(in) begin
		sadas
	end

endmodule 