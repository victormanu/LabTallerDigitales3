module ALU(in,out);
	input logic in;
	input logic out;
	
	always @(in) begin
		in = in + 1;
	end

endmodule 