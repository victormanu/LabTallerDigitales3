module multiplicacion(a,b,c);
	input logic a;
	input logic b;
	output logic c;
endmodule
