module ALU();


endmodule 